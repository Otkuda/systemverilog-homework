//----------------------------------------------------------------------------
// Example
//----------------------------------------------------------------------------

module sort_two_floats_ab (
    input        [FLEN - 1:0] a,
    input        [FLEN - 1:0] b,

    output logic [FLEN - 1:0] res0,
    output logic [FLEN - 1:0] res1,
    output                    err
);

    logic a_less_or_equal_b;

    f_less_or_equal i_floe (
        .a   ( a                 ),
        .b   ( b                 ),
        .res ( a_less_or_equal_b ),
        .err ( err               )
    );

    always_comb begin : a_b_compare
        if ( a_less_or_equal_b ) begin
            res0 = a;
            res1 = b;
        end
        else
        begin
            res0 = b;
            res1 = a;
        end
    end

endmodule

//----------------------------------------------------------------------------
// Example - different style
//----------------------------------------------------------------------------

module sort_two_floats_array
(
    input        [0:1][FLEN - 1:0] unsorted,
    output logic [0:1][FLEN - 1:0] sorted,
    output                         err
);

    logic u0_less_or_equal_u1;

    f_less_or_equal i_floe
    (
        .a   ( unsorted [0]        ),
        .b   ( unsorted [1]        ),
        .res ( u0_less_or_equal_u1 ),
        .err ( err                 )
    );

    always_comb
        if (u0_less_or_equal_u1)
            sorted = unsorted;
        else
              {   sorted [0],   sorted [1] }
            = { unsorted [1], unsorted [0] };

endmodule

//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module sort_three_floats (
    input        [0:2][FLEN - 1:0] unsorted,
    output logic [0:2][FLEN - 1:0] sorted,
    output                         err
);

    // Task:
    // Implement a module that accepts three Floating-Point numbers and outputs them in the increasing order.
    // The module should be combinational with zero latency.
    // The solution can use up to three instances of the "f_less_or_equal" module.
    //
    // Notes:
    // res0 must be less or equal to the res1
    // res1 must be less or equal to the res2
    //
    // The FLEN parameter is defined in the "import/preprocessed/cvw/config-shared.vh" file
    // and usually equal to the bit width of the double-precision floating-point number, FP64, 64 bits.
    logic f0_leq_f1, f1_leq_f2;
    logic err1, err2, err3;
    // temps for preventing loopbacks in comb logic
    logic [0:1][FLEN-1:0] presorted; // temporary result after 1st comp
    logic [FLEN-1:0] presorted_1;   // temporary result after 2 comp


    f_less_or_equal i_floe_0
    (
        .a   ( unsorted [0] ),
        .b   ( unsorted [1] ),
        .res ( f0_leq_f1    ),
        .err ( err1         )
    );

    f_less_or_equal i_floe_1
    (
        .a   ( presorted [1] ),
        .b   ( unsorted  [2] ),
        .res ( f1_leq_f2    ),
        .err ( err2         )
    );

    f_less_or_equal i_floe_2
    (
        .a   ( presorted [0] ),
        .b   ( presorted_1 ),
        .res ( f0_leq_f1_s  ),
        .err ( err3         )
    );


    always_comb begin
      if (!f0_leq_f1) { presorted[0], presorted[1] } = { unsorted[1], unsorted[0] };
      else presorted[0:1] = unsorted[0:1];

      if (!f1_leq_f2) { presorted_1, sorted[2] } = { unsorted[2], presorted[1] };
      else { presorted_1, sorted[2] } = { presorted[1], unsorted[2] };

      if (!f0_leq_f1_s) {sorted[0], sorted[1]} = { presorted_1, presorted[0] };
      else {sorted[0], sorted[1]} = { presorted[0], presorted_1 };
    end

    assign err = err1 | err2 | err3;


endmodule
